// Writeback Stage
module writeback (
    // ports
);
    
endmodule
