module Clk_generator(clk);
    output reg clk;

    
endmodule