`ifndef BUTTONS
`define BUTTONS

module buttons(
    input clk, //Main clk
    output [1:0] buttons_output //The output from the buttons
);

    

endmodule

`endif