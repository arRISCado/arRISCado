// Execute Stage
module execute (
    // ports
);
    
endmodule
