`ifndef BUTTONS
`define BUTTONS

module buttons(
    input clk, //Main clk
    input btn1,
    input btn2,
    output [1:0] buttons_output //The output from the buttons
);



endmodule

`endif