// Top Level Target for Primer 20k
module primer20k (
    // ports
);
    
endmodule
