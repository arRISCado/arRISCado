// Memory Stage
module memory (
    // ports
);
    
endmodule
