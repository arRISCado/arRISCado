// Decode Stage
module decode (
    // ports
);
    
endmodule
