// Memory Management Unit
module mmu (
    // ports
);
    
endmodule
