module top(clk);
    input clk;

    Processor processor(clk);

endmodule