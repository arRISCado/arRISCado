// Top Level Target for Primer 20k
`include "../../project/cpu.v"

module primer20k (
    // ports
);
    
endmodule
