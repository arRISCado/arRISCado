// Arithmetic Logic Unit
module alu (
  // ports
);

endmodule
