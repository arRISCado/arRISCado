module Memory(clk, addr, w_data, r_data, w_enable, r_enable);
    input [31:0] addr, w_data;
    output r_data;
    input w_enable, r_enable;

endmodule