// Fetch Stage
module fetch (
    // ports
);
    
endmodule
