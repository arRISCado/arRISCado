// Top Level Target for Nano 20k
module nano20k (
    // ports
);
    
endmodule
